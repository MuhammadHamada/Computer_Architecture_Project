LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;

ENTITY ROM IS  
	PORT ( 
		data    :   OUT STD_LOGIC_VECTOR(24 downto 0);
		ADDRESS :   IN  STD_LOGIC_VECTOR (4 DOWNTO 0) 
		);    
END ENTITY ROM;


ARCHITECTURE DATAFLOW  OF ROM IS

TYPE ROM_TYPE IS ARRAY(0 TO 31) of std_logic_vector(24 DOWNTO 0);
     SIGNAL ROM : ROM_TYPE :=(
   0     => "1100100010101110000000001",
   1     => "0010001100110000001000000",
   2     => "1101000110011110110001000",
   3     => "1100010011001110000000101",
   4     => "1101001000011111110001000",
   5     => "0010001100100000000000000",
   6     => "1100100010101110000000111",
   7     => "0011000000001111110001000",
   8     => "0001111011110000000000000",
   9     => "1100111111010000010001000",
   10    => "1001010111101110100001000",
   11    => "1100100010101110000010001",
   12    => "1101011001101111100001000",
   13    => "0001111010000000000000000",
   14    => "1100100010101110000001111",
   15    => "0011010000000011100001000",
   16    => "0100001101100000000000000",
   17    => "1100111111010000000010011",
   18    => "0101010111100110000100000",
   19    => "1000010101000111000111001",
   20    => "0101011001100111000100000",
   21    => "1010110000000011000011111",
   22    => "1100100010101110000010101",
   23    => "1100010010101110000010101",
   24    => "0010001101100000000000000",
   25    => "0110001100100000000000000",
   26    => "1101010111100010000100000",
   27    => "1100001110000000000000000",
   28    =>  "1101011001100011000100000",
   29    => "1110100000100000000000000",
   30    => "1100111111010000000010111",
   31    => "0000001100001000000100000"
);

BEGIN

data <= ROM(to_integer(unsigned(ADDRESS))) ;

END DATAFLOW;